----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 09/22/2025 09:18:19 PM
-- Design Name: Eyosiyas Endalamaw
-- Module Name: decoder - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity decoder is
  Port (
  clk : in std_logic;
  --reset : in std_logic;
  eyu : in std_logic_vector(31 downto 0); -- this one is used for accepting the insert values.
  Asel : out std_logic_vector(4 downto 0);
  Bsel : out std_logic_vector(4 downto 0);
  Dsel : out std_logic_vector(4 downto 0);
  Dlen : out std_logic;
  PCAsel : out std_logic;
  IMMBsel : out std_logic;
  IMM : out std_logic_vector(31 downto 0);
  PCDsel : out std_logic;
  PCle : out std_logic;
  PCie : out std_logic;
  isBr : out std_logic;
  BRcond : out std_logic_vector(2 downto 0);
  ALUfunc : out std_logic_vector(3 downto 0);
  eyu_illegal : out std_logic  --- this one is used to catch illegal values.
   );
end decoder;

architecture Behavioral of decoder is

     -- opcode constants 
     constant OPC_OP : std_logic_vector(6 downto 0) := "0110011"; -- R-type
     constant OPC_OPIMM : std_logic_vector(6 downto 0) := "0010011"; -- I-type ALU
     constant OPC_load : std_logic_vector(6 downto 0) := "0000011"; -- Load
     constant OPC_store : std_logic_vector(6 downto 0) := "0100011"; -- store
     constant OPC_branch : std_logic_vector(6 downto 0) := "1100011"; -- branches
     constant OPC_JALR : std_logic_vector(6 downto 0) := "1100111"; -- JALR
     constant OPC_JAL : std_logic_vector(6 downto 0) := "1101111"; -- JAL
     constant OPC_lui : std_logic_vector(6 downto 0) := "0110111"; -- LUI
     constant OPC_AUIPC : std_logic_vector(6 downto 0) := "0010111"; -- AUIPC
     constant OPC_System : std_logic_vector(6 downto 0) := "1110011"; -- system (ecall/ebreak/csr)
     constant OPC_MISC : std_logic_vector(6 downto 0) := "0001111"; -- Fench
     
     -- alu function constants 
     constant ALU_add : std_logic_vector (3 downto 0) := "0000";
     constant ALU_sub : std_logic_vector (3 downto 0) := "0001";
     constant ALU_and : std_logic_vector (3 downto 0) := "0010";
     constant ALU_or : std_logic_vector (3 downto 0) := "0011";
     constant ALU_xor : std_logic_vector (3 downto 0) := "0100";
     constant ALU_slt : std_logic_vector (3 downto 0) := "0101";
     constant ALU_sltu : std_logic_vector (3 downto 0) := "0110";
     constant ALU_sll : std_logic_vector (3 downto 0) := "0111";
     constant ALU_srl : std_logic_vector (3 downto 0) := "1000";
     constant ALU_sra : std_logic_vector (3 downto 0) := "1001";
     
     -- extract fields from the table imm (funct7), rs2, rs2, funct3, rd, opcode
     signal opcode : std_logic_vector(6 downto 0);
     signal rd : std_logic_vector(4 downto 0);
     signal funct3 : std_logic_vector(2 downto 0);
     signal rs1 : std_logic_vector(4 downto 0);
     signal rs2 : std_logic_vector(4 downto 0);
     signal funct7 : std_logic_vector(6 downto 0);
     
     -- extend the bits into 32bit 
     function set_extend32(x : std_logic_vector) return std_logic_vector is 
     begin
         return std_logic_vector(RESIZE(signed(x), 32));
     end;
     
     -- extract the immediate values from the 32-bit.
     --for I-type
     function imm_i(eyu : std_logic_vector(31 downto 0)) return std_logic_vector is
     variable raw : std_logic_vector(11 downto 0);
     begin
          raw := eyu(31 downto 20);
          return set_extend32(raw);
     end;
     
     -- for S-type 
     function imm_s(eyu : std_logic_vector(31 downto 0)) return std_logic_vector is
     variable raw : std_logic_vector(11 downto 0);
     begin
          raw := eyu(31 downto 25) & eyu(11 downto 7);
          return set_extend32(raw);
     end;
     
     --for B-type
     function imm_b(eyu : std_logic_vector(31 downto 0)) return std_logic_vector is
     variable raw : std_logic_vector(12 downto 0);
     begin
          raw := eyu(31) & eyu(7) & eyu(30 downto 25) & eyu(11 downto 8) & '0';
          return set_extend32(raw);
     end;
     
     -- for U type
     function imm_u(eyu : std_logic_vector(31 downto 0)) return std_logic_vector is
     begin
          return eyu(31 downto 12) & (11 downto 0 => '0');
     end;
     
     -- J-type
     function imm_j(eyu : std_logic_vector(31 downto 0)) return std_logic_vector is
     variable raw : std_logic_vector(20 downto 0);
     begin
          raw := eyu(31) & eyu(19 downto 12) & eyu(20) & eyu(30 downto 21) & '0';
          return set_extend32(raw);
     end;
     
     -- translate funct3 into branch BRcond
     function map_brcond(f3 : std_logic_vector(2 downto 0)) return std_logic_vector is
     begin
        case f3 is 
            when "000" => return "000"; --BEQ
            when "001" => return "001"; --BNEQ
            when "010" => return "010"; --BLT
            when "011" => return "011"; --BGE
            when "110" => return "110"; --BLTU
            when "111" => return "111"; --BGEU
            when others => return "000";
        end case;
     end;
     
     -- Decode ALU function for op and op-imm
     function decoder_alu(opcode : std_logic_vector(6 downto 0);
                          f3 : std_logic_vector(2 downto 0);
                          f7 : std_logic_vector(6 downto 0))
                          return std_logic_vector  is
     begin
         if opcode = OPC_OP then
            case f3 is
                when "000" => if f7 = "0100000" then return ALU_SUB; else return ALU_ADD; end if;
                when "001" => return ALU_sll;
                when "010" => return ALU_slt;
                when "011" => return ALU_sltu;
                when "100" => return ALU_xor;
                when "101" => if f7 = "0100000" then return ALU_sra; else return ALU_srl; end if;
                when "110" => return ALU_or;
                when "111" => return ALU_and;
                when others => return ALU_add;
            end case;
         elsif opcode = OPC_OPIMM then
            case f3 is
               when "000" => return ALU_add; --addi
               when "010" => return ALU_slt;
               when "011" => return ALU_sltu;
               when "100" => return ALU_xor;
               when "110" => return ALU_or;
               when "111" => return ALU_and;
               when "001" => return ALU_sll;
               when "101" => if f7 = "0100000" then return ALU_sra; else return ALU_srl; end if;
               when others => return ALU_add;
            end case;
         else
             return ALU_add;
         end if;
     
     end;

begin

    -- field extraction sections
    opcode <= eyu(6 downto 0);
    rd <= eyu(11 downto 7);
    funct3 <= eyu(14 downto 12);
    rs1 <= eyu(19 downto 15);
    rs2 <= eyu(24 downto 20);
    funct7 <= eyu(31 downto 25);
    
    process(opcode, rs1, rs2, rd, funct3, funct7, eyu)
        -- tempo variable storage
        variable v_Asel : std_logic_vector(4 downto 0) := (others => '0');
        variable v_Bsel : std_logic_vector(4 downto 0) := (others => '0');
        variable v_Dsel : std_logic_vector(4 downto 0) := (others => '0');
        variable v_Dlen : std_logic := '0';
        variable v_PCAsel : std_logic := '0';
        variable v_IMMBsel : std_logic := '0';
        variable v_IMM : std_logic_vector(31 downto 0) := (others => '0');
        variable v_PCDsel : std_logic := '0';
        variable v_PCle : std_logic := '0';
        variable v_PCie : std_logic := '0';
        variable v_isBr : std_logic := '0';
        variable v_BRcond : std_logic_vector(2 downto 0) := "000";
        variable v_ALUfunc : std_logic_vector(3 downto 0) := ALU_add;
        variable v_eyu_illegal : std_logic := '0';
            
    begin
        -- passing rs1, rs2, rd into v_Asel, v_Bsel, v_Dsel
        v_Asel := rs1;
        v_Bsel := rs2;
        v_Dsel := rd;
        
        case opcode is
            -- R-type ALU
            when OPC_OP =>
                v_Dlen := '1';
                v_IMMBsel := '0'; --rs2
                v_PCAsel := '0';
                v_PCDsel := '0';
                v_ALUfunc := decoder_alu(opcode, funct3, funct7);
                v_eyu_illegal := '0';
                
             -- I-type ALU
            when OPC_OPIMM =>
                v_Dlen := '1';
                v_IMMBsel := '1'; --imm
                v_PCAsel := '0';
                v_PCDsel := '0';
                v_IMM := imm_i(eyu);
                v_ALUfunc := decoder_alu(opcode, funct3, funct7);
                v_eyu_illegal := '0';
                
            -- load
            when OPC_load =>
                v_Dlen := '0';
                v_IMMBsel := '1';
                v_PCAsel := '0';
                v_PCDsel := '0';
                v_IMM := imm_i(eyu);
                v_ALUfunc := ALU_add;
                v_eyu_illegal := '0';
                
             -- store
            when OPC_store =>
                v_Dlen := '0';
                v_IMMBsel := '1';
                v_PCAsel := '0';
                v_PCDsel := '0';
                v_IMM := imm_s(eyu);
                v_ALUfunc := ALU_add;
                v_eyu_illegal := '0';
                
             -- branches
            when OPC_branch =>
                v_Dlen := '0';
                v_IMMBsel := '1';
                v_PCAsel := '1';
                v_PCDsel := '0';
                v_IMM := imm_b(eyu);
                v_ALUfunc := ALU_add;
                v_isBR := '1';
                v_BRcond := map_brcond(funct3);
                v_PCle := '0';
                v_eyu_illegal := '0';
                
            -- jal
            when OPC_JAL =>
                v_isBR := '0';
                v_IMMBsel := '1';
                v_PCAsel := '1';
                v_IMM := imm_j(eyu);
                v_ALUfunc := ALU_add;
                v_PCle := '1';
                v_Dlen := '0';
                v_eyu_illegal := '0';
                
             -- jalr
            when OPC_JALR =>
                v_IMMBsel := '1';
                v_PCAsel := '0';
                v_IMM := imm_i(eyu);
                v_ALUfunc := ALU_add;
                v_PCle := '1';
                v_Dlen := '0';
                v_eyu_illegal := '0';
                
            -- lui
            when OPC_lui =>
                v_Asel := "00000";
                v_IMMBsel := '1';
                v_PCAsel := '0';
                v_PCDsel := '0';
                v_IMM := imm_u(eyu);
                v_ALUfunc := ALU_add;
                v_Dlen := '1';
                v_eyu_illegal := '0';
                
            -- auipc
            when OPC_AUIPC =>
                v_PCAsel := '1';
                v_IMMBsel := '1';
                v_PCDsel := '0';
                v_ALUfunc := ALU_add;
                v_Dlen := '1';
                v_IMM := imm_u(eyu);    
                v_eyu_illegal := '0';
                
            -- stystem 
            when OPC_System | OPC_MISC =>
                 v_Dlen := '0';    
                
            when others => v_eyu_illegal := '1';  
        
        end case;
        
        --move this tempo values into the outputs
        Asel <= v_Asel;
        Bsel <= v_Bsel;
        Dsel <= v_Dsel;
        Dlen <= v_Dlen;
        PCAsel <= v_PCAsel;
        IMMBsel <= v_IMMBsel;
        PCDsel <= v_PCDsel;
        PCle <= v_PCle;
        PCie <= v_PCie;
        isBR <= v_isBR;
        BRcond <= v_BRcond;
        ALUfunc <= v_ALUfunc;
        IMM <= v_IMM;
        eyu_illegal <= v_eyu_illegal;
        
    end process;

end Behavioral;








































