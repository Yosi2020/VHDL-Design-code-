----------------------------------------------------------------------------------
-- Company: sdsmt
-- Engineer: Eyosiyas
-- 
-- Create Date: 09/02/2025 11:33:10 AM
-- Design Name: Eyosiyas
-- Module Name: lab1 - Behavioral
-- Project Name: Lab1 ALUFUNC
-- Target Devices: None
-- Tool Versions: v1.0
-- Description: None
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity data_path is
  Port ( 
  clk : in std_logic;
  reset : in std_logic;
  Asel : in std_logic_vector(4 downto 0);
  Bsel : in std_logic_vector(4 downto 0);
  Dsel : in std_logic_vector(4 downto 0);
  Dlen : in std_logic;
  PCAsel : in std_logic;
  IMMBsel : in std_logic;
  PCDsel : in std_logic;
  PCle : in std_logic;
  PCie : in std_logic;
  isBR : in std_logic;
  BRcond : std_logic_vector(2 downto 0);
  ALUFunc : std_logic_vector(3 downto 0);
  IMM : std_logic_vector(31 downto 0);
  PC_q : out std_logic_vector(31 downto 0);
  alu_y : out std_logic_vector(31 downto 0);
  regA_q : out std_logic_vector(31 downto 0);
  regB_q : out std_logic_vector(31 downto 0)
  --branch_q : out std_logic
  );
end data_path;

architecture Behavioral of data_path is
    signal Abus, Bbus : std_logic_vector(31 downto 0);
    signal Dbus : std_logic_vector(31 downto 0);
    signal RegA : std_logic_vector(31 downto 0);
    signal RegB : std_logic_vector(31 downto 0);
    signal ALU_out : std_logic_vector(31 downto 0);
    signal pc_out : std_logic_vector(31 downto 0);
    signal PCle_sig : std_logic;
     
begin
    U_REG : entity work.regsiter_file port map 
    (
    clk => clk,
    reset => reset,
    Asel => Asel,
    Bsel => Bsel,
    Dsel => Dsel,
    Dlen => Dlen,
    Dbus => Dbus,
    Aout => RegA,
    Bout => RegB
    );
    
    
    regA_q <= RegA;
    regB_q <= RegB;
    
    U_ALU : entity work.alu port map (
    clk => clk,
    reset => reset,
    Aout => REGA,
    Bout => REGB,
    PCAsel => PCAsel,
    IMM => IMM,
    IMMBsel => IMMBsel,
    PCout => pc_out,
    ALUfun => ALUFunc,
    eyu_out => ALU_out
    );
    
    alu_y <= ALU_out;
    
    U_BRANCH : entity work.branch port map (
    clk => clk,
    reset => reset,
    isBR => isBR,
    BRcond => BRcond,
    A => REGA,
    B => REGB,
    eyu_output => PCle_sig
    );
    
    --branch_q <= PCle_sig;
    
    U_PC : entity work.PC port map(
    clk => clk,
    reset => reset,
    PCle => PCle,
    PCie => PCie,
    Branch_out => PCle_sig,
    ALUout => ALU_out,
    eyu_out => pc_out
    );
    
    pc_q <= pc_out;
    
    Dbus <= PC_out when PCDsel = '1' else ALU_out;
    
   
end Behavioral;
